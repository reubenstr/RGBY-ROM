// Convert 8-bit value into sinusoid equivalent.
// Generated from generateSin.py

module sinTable(
input [7:0] in,
output [7:0] out);

assign out =
	(in == 0) ? 0 :
	(in == 1) ? 0 :
	(in == 2) ? 0 :
	(in == 3) ? 0 :
	(in == 4) ? 0 :
	(in == 5) ? 0 :
	(in == 6) ? 0 :
	(in == 7) ? 0 :
	(in == 8) ? 1 :
	(in == 9) ? 1 :
	(in == 10) ? 1 :
	(in == 11) ? 1 :
	(in == 12) ? 1 :
	(in == 13) ? 2 :
	(in == 14) ? 2 :
	(in == 15) ? 2 :
	(in == 16) ? 2 :
	(in == 17) ? 3 :
	(in == 18) ? 3 :
	(in == 19) ? 3 :
	(in == 20) ? 4 :
	(in == 21) ? 4 :
	(in == 22) ? 5 :
	(in == 23) ? 5 :
	(in == 24) ? 5 :
	(in == 25) ? 6 :
	(in == 26) ? 6 :
	(in == 27) ? 7 :
	(in == 28) ? 7 :
	(in == 29) ? 8 :
	(in == 30) ? 9 :
	(in == 31) ? 9 :
	(in == 32) ? 10 :
	(in == 33) ? 10 :
	(in == 34) ? 11 :
	(in == 35) ? 12 :
	(in == 36) ? 12 :
	(in == 37) ? 13 :
	(in == 38) ? 14 :
	(in == 39) ? 14 :
	(in == 40) ? 15 :
	(in == 41) ? 16 :
	(in == 42) ? 17 :
	(in == 43) ? 17 :
	(in == 44) ? 18 :
	(in == 45) ? 19 :
	(in == 46) ? 20 :
	(in == 47) ? 21 :
	(in == 48) ? 21 :
	(in == 49) ? 22 :
	(in == 50) ? 23 :
	(in == 51) ? 24 :
	(in == 52) ? 25 :
	(in == 53) ? 26 :
	(in == 54) ? 27 :
	(in == 55) ? 28 :
	(in == 56) ? 29 :
	(in == 57) ? 30 :
	(in == 58) ? 31 :
	(in == 59) ? 32 :
	(in == 60) ? 33 :
	(in == 61) ? 34 :
	(in == 62) ? 35 :
	(in == 63) ? 36 :
	(in == 64) ? 37 :
	(in == 65) ? 38 :
	(in == 66) ? 40 :
	(in == 67) ? 41 :
	(in == 68) ? 42 :
	(in == 69) ? 43 :
	(in == 70) ? 44 :
	(in == 71) ? 45 :
	(in == 72) ? 47 :
	(in == 73) ? 48 :
	(in == 74) ? 49 :
	(in == 75) ? 50 :
	(in == 76) ? 52 :
	(in == 77) ? 53 :
	(in == 78) ? 54 :
	(in == 79) ? 55 :
	(in == 80) ? 57 :
	(in == 81) ? 58 :
	(in == 82) ? 59 :
	(in == 83) ? 61 :
	(in == 84) ? 62 :
	(in == 85) ? 63 :
	(in == 86) ? 65 :
	(in == 87) ? 66 :
	(in == 88) ? 67 :
	(in == 89) ? 69 :
	(in == 90) ? 70 :
	(in == 91) ? 72 :
	(in == 92) ? 73 :
	(in == 93) ? 74 :
	(in == 94) ? 76 :
	(in == 95) ? 77 :
	(in == 96) ? 79 :
	(in == 97) ? 80 :
	(in == 98) ? 82 :
	(in == 99) ? 83 :
	(in == 100) ? 85 :
	(in == 101) ? 86 :
	(in == 102) ? 88 :
	(in == 103) ? 89 :
	(in == 104) ? 90 :
	(in == 105) ? 92 :
	(in == 106) ? 93 :
	(in == 107) ? 95 :
	(in == 108) ? 97 :
	(in == 109) ? 98 :
	(in == 110) ? 100 :
	(in == 111) ? 101 :
	(in == 112) ? 103 :
	(in == 113) ? 104 :
	(in == 114) ? 106 :
	(in == 115) ? 107 :
	(in == 116) ? 109 :
	(in == 117) ? 110 :
	(in == 118) ? 112 :
	(in == 119) ? 113 :
	(in == 120) ? 115 :
	(in == 121) ? 117 :
	(in == 122) ? 118 :
	(in == 123) ? 120 :
	(in == 124) ? 121 :
	(in == 125) ? 123 :
	(in == 126) ? 124 :
	(in == 127) ? 126 :
	(in == 128) ? 128 :
	(in == 129) ? 129 :
	(in == 130) ? 131 :
	(in == 131) ? 132 :
	(in == 132) ? 134 :
	(in == 133) ? 135 :
	(in == 134) ? 137 :
	(in == 135) ? 138 :
	(in == 136) ? 140 :
	(in == 137) ? 142 :
	(in == 138) ? 143 :
	(in == 139) ? 145 :
	(in == 140) ? 146 :
	(in == 141) ? 148 :
	(in == 142) ? 149 :
	(in == 143) ? 151 :
	(in == 144) ? 152 :
	(in == 145) ? 154 :
	(in == 146) ? 155 :
	(in == 147) ? 157 :
	(in == 148) ? 158 :
	(in == 149) ? 160 :
	(in == 150) ? 162 :
	(in == 151) ? 163 :
	(in == 152) ? 165 :
	(in == 153) ? 166 :
	(in == 154) ? 167 :
	(in == 155) ? 169 :
	(in == 156) ? 170 :
	(in == 157) ? 172 :
	(in == 158) ? 173 :
	(in == 159) ? 175 :
	(in == 160) ? 176 :
	(in == 161) ? 178 :
	(in == 162) ? 179 :
	(in == 163) ? 181 :
	(in == 164) ? 182 :
	(in == 165) ? 183 :
	(in == 166) ? 185 :
	(in == 167) ? 186 :
	(in == 168) ? 188 :
	(in == 169) ? 189 :
	(in == 170) ? 190 :
	(in == 171) ? 192 :
	(in == 172) ? 193 :
	(in == 173) ? 194 :
	(in == 174) ? 196 :
	(in == 175) ? 197 :
	(in == 176) ? 198 :
	(in == 177) ? 200 :
	(in == 178) ? 201 :
	(in == 179) ? 202 :
	(in == 180) ? 203 :
	(in == 181) ? 205 :
	(in == 182) ? 206 :
	(in == 183) ? 207 :
	(in == 184) ? 208 :
	(in == 185) ? 210 :
	(in == 186) ? 211 :
	(in == 187) ? 212 :
	(in == 188) ? 213 :
	(in == 189) ? 214 :
	(in == 190) ? 215 :
	(in == 191) ? 217 :
	(in == 192) ? 218 :
	(in == 193) ? 219 :
	(in == 194) ? 220 :
	(in == 195) ? 221 :
	(in == 196) ? 222 :
	(in == 197) ? 223 :
	(in == 198) ? 224 :
	(in == 199) ? 225 :
	(in == 200) ? 226 :
	(in == 201) ? 227 :
	(in == 202) ? 228 :
	(in == 203) ? 229 :
	(in == 204) ? 230 :
	(in == 205) ? 231 :
	(in == 206) ? 232 :
	(in == 207) ? 233 :
	(in == 208) ? 234 :
	(in == 209) ? 234 :
	(in == 210) ? 235 :
	(in == 211) ? 236 :
	(in == 212) ? 237 :
	(in == 213) ? 238 :
	(in == 214) ? 238 :
	(in == 215) ? 239 :
	(in == 216) ? 240 :
	(in == 217) ? 241 :
	(in == 218) ? 241 :
	(in == 219) ? 242 :
	(in == 220) ? 243 :
	(in == 221) ? 243 :
	(in == 222) ? 244 :
	(in == 223) ? 245 :
	(in == 224) ? 245 :
	(in == 225) ? 246 :
	(in == 226) ? 246 :
	(in == 227) ? 247 :
	(in == 228) ? 248 :
	(in == 229) ? 248 :
	(in == 230) ? 249 :
	(in == 231) ? 249 :
	(in == 232) ? 250 :
	(in == 233) ? 250 :
	(in == 234) ? 250 :
	(in == 235) ? 251 :
	(in == 236) ? 251 :
	(in == 237) ? 252 :
	(in == 238) ? 252 :
	(in == 239) ? 252 :
	(in == 240) ? 253 :
	(in == 241) ? 253 :
	(in == 242) ? 253 :
	(in == 243) ? 253 :
	(in == 244) ? 254 :
	(in == 245) ? 254 :
	(in == 246) ? 254 :
	(in == 247) ? 254 :
	(in == 248) ? 254 :
	(in == 249) ? 255 :
	(in == 250) ? 255 :
	(in == 251) ? 255 :
	(in == 252) ? 255 :
	(in == 253) ? 255 :
	(in == 254) ? 255 :
	(in == 255) ? 255 :
	0;
endmodule
